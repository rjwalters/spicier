RC Transient - Current Source Charging
I1 0 1 1m
R1 1 0 1k
C1 1 0 1u
.tran 10u 5m
.end
