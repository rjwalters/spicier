Voltage Divider with .PRINT
V1 1 0 10
R1 1 2 1k
R2 2 0 1k
.PRINT DC V(1) V(2)
.OP
.END
