Diode Circuit - R + D
V1 1 0 DC 5
R1 1 2 1k
D1 2 0
.op
.end
